  LIBRARY ieee;
  USE ieee.std_logic_1164.ALL;
  USE ieee.numeric_std.ALL;
  use work.ADAT.all;
  


  ENTITY tb_ADAT_Dekoder IS
  END tb_ADAT_Dekoder;

  ARCHITECTURE behavior OF tb_ADAT_Dekoder IS 
		constant SCHNITTSTELLEN : natural := 3;
		--#############################
  		signal tb_clk				: std_logic := '1';
  		signal tb_AdatIn        : bit;
		signal tb_AdatTakt      : std_logic;
		signal tb_AdatFramesync : std_logic := '0';
		------------------
  		signal tb_adat : bit_vector(0 to SCHNITTSTELLEN-1);
		signal tb_Out_Daten : ADAT_Daten_Array(0 to SCHNITTSTELLEN-1);
		signal tb_Out_FrameOK: bit_vector(0 to SCHNITTSTELLEN-1);
		
		COMPONENT ADAT_Taktgewinnung
		Port(clk 			  : in std_logic;
			  -- Daten-Eingang
			  In_ADAT 		  : in bit;
			  
			  -- Takt-Ausgang
			  Out_ADAT_Clock : out std_logic;
			  Frame_Sync     : out std_logic
			  );
		END COMPONENT;
		
		COMPONENT ADAT_Dekoder
		generic (AdatSchnittstellen : integer := 3);
		Port(ADAT_Takt		  : in std_logic;
			  ADAT_Sync		  : in bit;
			  -- Daten-Eing�nge
			  In_ADAT 		  : in bit_vector(0 to SCHNITTSTELLEN-1);
			  
			  -- Daten-Ausgang			  
			  Out_Daten 	  : out ADAT_Daten_Array(0 to AdatSchnittstellen-1);
			  Out_FrameOK    : out bit_vector(0 to AdatSchnittstellen-1);
			  Out_NeueDaten  : out bit
			  );
		END COMPONENT;
  BEGIN
		tb_clk  <= not tb_clk after 0.5 * 1.769134964 ns; --5ns -> 100MHz  
		----------[TAKT]-------------------------------------------------------------------------------------
		-- !!! TODO: L�sst sich entsch�rfen, weil das Sync-signal nicht relevant f�r die Daten ist !!!
		--
		-- Muss so gew�hlt werden, dass der Bitlaengenz�hler f�r einen Taktwechsel (halbe Periode)
		-- gr��er als 22 wird (10Bit+1Bit davor)*2Taktwechsel,
      --	damit auch im Sync die m�gliche Abweichung von 1Bit/Wechsel unter der Zeit f�r einen Takt bleibt.
		-- (wodurch sonst ein zus�tzlicher Wechsel in der ADAT-Taktleitung erzeugt werden w�rde)
		--
		-- Optimal: Periode = 1/(48000*2*256*23)
		--
		-- Sync:    	   _------------------------------------------------------------------_____
		-- Wechsel Nr: 	 01.02.03.04.05.06.07.08.09.10.11.12.13.14.15.16.17.18.19.20.21.22.
		-- Takt:          _---___---___---___---___---___---___---___---___---___---___---___---___
		-- Max. Abweichung:  1  2  3  4  5  6  7  8  9 10 11 12 13 14 15 16 17 18 19 20 21 22       
		--
		------------------------------------------------------------------------------------------------------
		
		
		
		
		--
		tb_adat(0) <= '1',
'0' after 49600 ps,
'1' after 130800 ps,
'0' after 214 ns,
'1' after 292 ns,
'0' after 376 ns,
'1' after 456 ns,
'0' after 539600 ps,
'1' after 617200 ps,
'0' after 700400 ps,
'1' after 781600 ps,
'0' after 864400 ps,
'1' after 943600 ps,
'0' after 1026400 ps,
'1' after 1106400 ps,
'0' after 1190400 ps,
'1' after 1268400 ps,
'0' after 1351600 ps,
'1' after 1432800 ps,
'0' after 1515600 ps,
'1' after 1594400 ps,
'0' after 1677600 ps,
'1' after 1839600 ps,
'0' after 1921600 ps,
'1' after 2002400 ps,
'0' after 2085200 ps,
'1' after 2164 ns,
'0' after 2246800 ps,
'1' after 2653200 ps,
'0' after 3061600 ps,
'1' after 3466 ns,
'0' after 3875200 ps,
'1' after 4279600 ps,
'0' after 4362400 ps,
'1' after 4688 ns,
'0' after 4769600 ps,
'1' after 4850400 ps,
'0' after 4933200 ps,
'1' after 5012 ns,
'0' after 5094800 ps,
'1' after 5175600 ps,
'0' after 5258800 ps,
'1' after 5337200 ps,
'0' after 5420800 ps,
'1' after 5501600 ps,
'0' after 5583600 ps,
'1' after 5663200 ps,
'0' after 5746 ns,
'1' after 5826400 ps,
'0' after 5909600 ps,
'1' after 5988400 ps,
'0' after 6070800 ps,
'1' after 6152400 ps,
'0' after 6234800 ps,
'1' after 6314400 ps,
'0' after 6396800 ps,
'1' after 6477600 ps,
'0' after 6560400 ps,
'1' after 6721200 ps,
'0' after 6803200 ps,
'1' after 6884800 ps,
'0' after 7130400 ps,
'1' after 7209200 ps,
'0' after 7292800 ps,
'1' after 7372400 ps,
'0' after 7456400 ps,
'1' after 7534 ns,
'0' after 7617600 ps,
'1' after 7698400 ps,
'0' after 7781200 ps,
'1' after 7860 ns,
'0' after 7943200 ps,
'1' after 8023600 ps,
'0' after 8106800 ps,
'1' after 8184800 ps,
'0' after 8268400 ps,
'1' after 8349600 ps,
'0' after 8432 ns,
'1' after 8511200 ps,
'0' after 8594400 ps,
'1' after 8674400 ps,
'0' after 8757600 ps,
'1' after 8836400 ps,
'0' after 8919600 ps,
'1' after 9162400 ps,
'0' after 9327200 ps,
'1' after 9569600 ps,
'0' after 9978400 ps,
'1' after 10382 ns,
'0' after 10791600 ps,
'1' after 11196400 ps,
'0' after 11442800 ps,
'1' after 11603600 ps,
'0' after 11850 ns,
'1' after 11928400 ps,
'0' after 12011200 ps,
'1' after 12091600 ps,
'0' after 12175200 ps,
'1' after 12253600 ps,
'0' after 12336800 ps,
'1' after 12417600 ps,
'0' after 12500800 ps,
'1' after 12579200 ps,
'0' after 12662400 ps,
'1' after 12743200 ps,
'0' after 12826 ns,
'1' after 12905200 ps,
'0' after 12988400 ps,
'1' after 13068400 ps,
'0' after 13152 ns,
'1' after 13230400 ps,
'0' after 13313200 ps,
'1' after 13394 ns,
'0' after 13477200 ps,
'1' after 13556 ns,
'0' after 13638800 ps,
'1' after 13719200 ps,
'0' after 13802800 ps,
'1' after 13881200 ps,
'0' after 14046800 ps,
'1' after 14126 ns,
'0' after 14209200 ps,
'1' after 14288400 ps,
'0' after 14371200 ps,
'1' after 14452 ns,
'0' after 15349200 ps,
'1' after 15753600 ps,
'0' after 16163200 ps,
'1' after 16567600 ps,
'0' after 16977200 ps,
'1' after 17381200 ps,
'0' after 17546400 ps,
'1' after 17707600 ps,
'0' after 17789200 ps,
'1' after 18114800 ps,
'0' after 18196400 ps,
'1' after 18277200 ps,
'0' after 18360400 ps,
'1' after 18439200 ps,
'0' after 18522 ns,
'1' after 18602800 ps,
'0' after 18686400 ps,
'1' after 18764800 ps,
'0' after 18848 ns,
'1' after 18928 ns,
'0' after 19011600 ps,
'1' after 19090 ns,
'0' after 19173200 ps,
'1' after 19253600 ps,
'0' after 19336800 ps,
'1' after 19415600 ps,
'0' after 19498800 ps,
'1' after 19578800 ps,
'0' after 19662800 ps,
'1' after 19741200 ps,
'0' after 19824 ns,
'1' after 19904800 ps,
'0' after 19987600 ps,
'1' after 20066800 ps,
'0' after 20149600 ps,
'1' after 20230800 ps,
'0' after 20476 ns,
'1' after 20555200 ps,
'0' after 20638800 ps,
'1' after 20718 ns,
'0' after 20802400 ps,
'1' after 20880 ns,
'0' after 20963200 ps,
'1' after 21044 ns,
'0' after 21127200 ps,
'1' after 21205600 ps,
'0' after 21289200 ps,
'1' after 21368800 ps,
'0' after 21452800 ps,
'1' after 21530400 ps,
'0' after 21614400 ps,
'1' after 21695200 ps,
'0' after 21778 ns,
'1' after 21856800 ps,
'0' after 21940400 ps,
'1' after 22020800 ps,
'0' after 22103600 ps,
'1' after 22182 ns,
'0' after 22265600 ps,
'1' after 22346 ns,
'0' after 22428800 ps,
'1' after 22670800 ps,
'0' after 22917200 ps,
'1' after 23078 ns,
'0' after 23160400 ps,
'1' after 23241200 ps,
'0' after 23324 ns,
'1' after 23402400 ps,
'0' after 23486 ns,
'1' after 23566800 ps,
'0' after 23650 ns,
'1' after 23727200 ps,
'0' after 23811200 ps,
'1' after 23892 ns,
'0' after 23975200 ps,
'1' after 24053600 ps,
'0' after 24136400 ps,
'1' after 24217600 ps,
'0' after 24300400 ps,
'1' after 24379200 ps,
'0' after 24462 ns,
'1' after 24542800 ps,
'0' after 24626 ns,
'1' after 24705200 ps,
'0' after 24787600 ps,
'1' after 24868400 ps,
'0' after 24951600 ps,
'1' after 25112 ns,
'0' after 25276400 ps,
'1' after 25438400 ps,
'0' after 25520400 ps,
'1' after 25600800 ps,
'0' after 25684 ns,
'1' after 25762 ns,
'0' after 25845600 ps,
'1' after 25926400 ps,
'0' after 26009200 ps,
'1' after 26088 ns,
'0' after 26170800 ps,
'1' after 26252 ns,
'0' after 26334800 ps,
'1' after 26413600 ps,
'0' after 26496400 ps,
'1' after 26577600 ps,
'0' after 26660 ns,
'1' after 26738800 ps,
'0' after 26822400 ps,
'1' after 26902800 ps,
'0' after 26986 ns,
'1' after 27064400 ps,
'0' after 27147600 ps,
'1' after 27228400 ps,
'0' after 27311200 ps,
'1' after 27472 ns,
'0' after 27554 ns,
'1' after 27717200 ps,
'0' after 27799600 ps,
'1' after 27960 ns,
'0' after 28042 ns,
'1' after 28123200 ps,
'0' after 28206400 ps,
'1' after 28285200 ps,
'0' after 28368 ns,
'1' after 28448800 ps,
'0' after 28531600 ps,
'1' after 28610800 ps,
'0' after 28693200 ps,
'1' after 28774 ns,
'0' after 28857200 ps,
'1' after 28936 ns,
'0' after 29018800 ps,
'1' after 29100 ns,
'0' after 29182800 ps,
'1' after 29261200 ps,
'0' after 29344 ns,
'1' after 29425200 ps,
'0' after 29508 ns,
'1' after 29587200 ps,
'0' after 29670 ns,
'1' after 29750400 ps,
'0' after 29914800 ps,
'1' after 29994 ns,
'0' after 30078 ns,
'1' after 30319600 ps,
'0' after 30402400 ps,
'1' after 30483600 ps,
'0' after 30565600 ps,
'1' after 30645200 ps,
'0' after 30728400 ps,
'1' after 30808 ns,
'0' after 30808400 ps,
'1' after 30808800 ps,
'0' after 30891600 ps,
'1' after 30970400 ps,
'0' after 31053600 ps,
'1' after 31134 ns,
'0' after 31217200 ps,
'1' after 31295600 ps,
'0' after 31378800 ps,
'1' after 31459600 ps,
'0' after 31542400 ps,
'1' after 31621200 ps,
'0' after 31704 ns,
'1' after 31784800 ps,
'0' after 31868 ns,
'1' after 31946800 ps,
'0' after 32030 ns,
'1' after 32110800 ps,
'0' after 32274800 ps,
'1' after 32354 ns,
'0' after 32437200 ps,
'1' after 32517200 ps,
'0' after 32682 ns,
'1' after 32842 ns,
'0' after 33251200 ps,
'1' after 33655600 ps,
'0' after 34065200 ps,
'1' after 34469600 ps,
'0' after 34797200 ps,
'1' after 34876400 ps,
'0' after 34959600 ps,
'1' after 35202800 ps,
'0' after 35284400 ps,
'1' after 36178 ns,
'0' after 36588400 ps,
'1' after 36992400 ps,
'0' after 37402 ns,
'1' after 37806 ns,
'0' after 38134400 ps,
'1' after 38214 ns,
'0' after 38541600 ps,
'1' after 38620 ns,
'0' after 38704 ns,
'1' after 38865200 ps,
'0' after 38947600 ps,
'1' after 39027600 ps,
'0' after 39111200 ps,
'1' after 39189600 ps,
'0' after 39272800 ps,
'1' after 39353200 ps,
'0' after 39436400 ps,
'1' after 39515200 ps,
'0' after 39598400 ps,
'1' after 39679200 ps,
'0' after 39762 ns,
'1' after 39841200 ps,
'0' after 39924 ns,
'1' after 40004400 ps,
'0' after 40087600 ps,
'1' after 40166400 ps,
'0' after 40249200 ps,
'1' after 40330400 ps,
'0' after 40412800 ps,
'1' after 40492 ns,
'0' after 40575200 ps,
'1' after 40655600 ps,
'0' after 40738800 ps,
'1' after 40980 ns,
'0' after 41062800 ps,
'1' after 41387600 ps,
'0' after 41469600 ps,
'1' after 41550400 ps,
'0' after 41550800 ps,
'1' after 41551200 ps,
'0' after 41633200 ps,
'1' after 41712800 ps,
'0' after 41796 ns,
'1' after 41875600 ps,
'0' after 41959200 ps,
'1' after 42037600 ps,
'0' after 42120800 ps,
'1' after 42202 ns,
'0' after 42284400 ps,
'1' after 42363200 ps,
'0' after 42446800 ps,
'1' after 42526800 ps,
'0' after 42610400 ps,
'1' after 42688 ns,
'0' after 42772 ns,
'1' after 42853200 ps,
'0' after 42935600 ps,
'1' after 43014400 ps,
'0' after 43097200 ps,
'1' after 43177600 ps,
'0' after 43261200 ps,
'1' after 43502800 ps,
'0' after 43830800 ps,
'1' after 43910 ns,
'0' after 44319200 ps,
'1' after 44722800 ps,
'0' after 45132400 ps,
'1' after 45536400 ps,
'0' after 45536800 ps,
'1' after 45537200 ps,
'0' after 45783200 ps,
'1' after 45944 ns,
'0' after 46353200 ps,
'1' after 46756800 ps,
'0' after 47166800 ps,
'1' after 47571200 ps,
'0' after 47981200 ps,
'1' after 48222 ns,
'0' after 48304800 ps,
'1' after 48386400 ps,
'0' after 48468400 ps,
'1' after 48791600 ps,
'0' after 48874 ns,
'1' after 48955200 ps,
'0' after 49038 ns,
'1' after 49116800 ps,
'0' after 49200 ns,
'1' after 49280400 ps,
'0' after 49364 ns,
'1' after 49442 ns,
'0' after 49525200 ps,
'1' after 49606800 ps,
'0' after 49689200 ps,
'1' after 49768 ns,
'0' after 49851200 ps,
'1' after 49931600 ps,
'0' after 50015200 ps,
'1' after 50093200 ps,
'0' after 50176400 ps,
'1' after 50257200 ps,
'0' after 50340400 ps,
'1' after 50418800 ps,
'0' after 50501600 ps,
'1' after 50582400 ps,
'0' after 50666 ns,
'1' after 50826400 ps,
'0' after 50908800 ps,
'1' after 50989600 ps,
'0' after 51072400 ps,
'1' after 51151600 ps,
'0' after 51234400 ps,
'1' after 51640400 ps,
'0' after 52049200 ps,
'1' after 52452800 ps,
'0' after 52863200 ps,
'1' after 53104400 ps,
'0' after 53269200 ps,
'1' after 53348400 ps,
'0' after 53514 ns,
'1' after 53674400 ps,
'0' after 54083600 ps,
'1' after 54487600 ps,
'0' after 54897200 ps,
'1' after 55301600 ps,
'0' after 55548 ns,
'1' after 55708800 ps,
'0' after 55873200 ps,
'1' after 55952800 ps,
'0' after 56036 ns,
'1' after 56115200 ps,
'0' after 57013600 ps,
'1' after 57417600 ps,
'0' after 57827600 ps,
'1' after 58232 ns,
'0' after 58641600 ps,
'1' after 59045200 ps,
'0' after 59210800 ps,
'1' after 59289600 ps,
'0' after 59455200 ps,
'1' after 59697200 ps,
'0' after 59861200 ps,
'1' after 59941600 ps,
'0' after 60025200 ps,
'1' after 60103200 ps,
'0' after 60186 ns,
'1' after 60266800 ps,
'0' after 60350400 ps,
'1' after 60428800 ps,
'0' after 60511600 ps,
'1' after 60593200 ps,
'0' after 60675600 ps,
'1' after 60754 ns,
'0' after 60837200 ps,
'1' after 60917600 ps,
'0' after 61001600 ps,
'1' after 61079200 ps,
'0' after 61162800 ps,
'1' after 61242800 ps,
'0' after 61327200 ps,
'1' after 61404800 ps,
'0' after 61488400 ps,
'1' after 61569200 ps,
'0' after 61733200 ps,
'1' after 61812 ns,
'0' after 61896 ns,
'1' after 62056800 ps,
'0' after 62303200 ps,
'1' after 62707200 ps,
'0' after 63116400 ps,
'1' after 63520800 ps,
'0' after 63930400 ps,
'1' after 64335200 ps,
'0' after 64743600 ps,
'1' after 65148 ns,
'0' after 65557600 ps,
'1' after 65962 ns,
'0' after 66371600 ps,
'1' after 66613200 ps,
'0' after 66777600 ps,
'1' after 66857600 ps,
'0' after 66941200 ps,
'1' after 67101200 ps,
'0' after 67184 ns,
'1' after 67590400 ps,
'0' after 67998400 ps,
'1' after 68402800 ps,
'0' after 68812800 ps,
'1' after 68891600 ps,
'0' after 68974800 ps,
'1' after 69217600 ps,
'0' after 69299200 ps,
'1' after 69380 ns,
'0' after 69463600 ps,
'1' after 69542400 ps,
'0' after 69625600 ps,
'1' after 70030400 ps,
'0' after 70440 ns,
'1' after 70844 ns,
'0' after 71253600 ps,
'1' after 71414400 ps,
'0' after 71660400 ps,
'1' after 71739600 ps,
'0' after 71823200 ps,
'1' after 71984 ns,
'0' after 72066 ns,
'1' after 72147200 ps,
'0' after 72230 ns,
'1' after 72308800 ps,
'0' after 72393200 ps,
'1' after 72471600 ps,
'0' after 72554800 ps,
'1' after 72635200 ps,
'0' after 72718400 ps,
'1' after 72797200 ps,
'0' after 72880 ns,
'1' after 72960800 ps,
'0' after 73044 ns,
'1' after 73122 ns,
'0' after 73205600 ps,
'1' after 73286 ns,
'0' after 73369200 ps,
'1' after 73448 ns,
'0' after 73530800 ps,
'1' after 73611600 ps,
'0' after 73694400 ps,
'1' after 73773200 ps,
'0' after 73938800 ps,
'1' after 74099600 ps,
'0' after 74264400 ps,
'1' after 74425200 ps,
'0' after 74507200 ps,
'1' after 74588400 ps,
'0' after 74671200 ps,
'1' after 74750 ns,
'0' after 74832800 ps,
'1' after 74913200 ps,
'0' after 74996800 ps,
'1' after 75075200 ps,
'0' after 75158 ns,
'1' after 75239200 ps,
'0' after 75322400 ps,
'1' after 75400400 ps,
'0' after 75484 ns,
'1' after 75564400 ps,
'0' after 75648400 ps,
'1' after 75726400 ps,
'0' after 75809200 ps,
'1' after 75890400 ps,
'0' after 75973200 ps,
'1' after 76052 ns,
'0' after 76135200 ps,
'1' after 76215200 ps,
'0' after 76299200 ps,
'1' after 76377200 ps,
'0' after 76542 ns,
'1' after 76622400 ps,
'0' after 76706 ns,
'1' after 76947600 ps,
'0' after 77845200 ps,
'1' after 78249600 ps,
'0' after 78332800 ps,
'1' after 78413600 ps,
'0' after 78496400 ps,
'1' after 78575600 ps,
'0' after 78659200 ps,
'1' after 78738400 ps,
'0' after 78822800 ps,
'1' after 78900800 ps,
'0' after 78984 ns,
'1' after 79064400 ps,
'0' after 79148 ns,
'1' after 79225600 ps,
'0' after 79309200 ps,
'1' after 79390800 ps,
'0' after 79472800 ps,
'1' after 79552 ns,
'0' after 79635200 ps,
'1' after 79714800 ps,
'0' after 79798800 ps,
'1' after 79876800 ps,
'0' after 79960800 ps,
'1' after 80041200 ps,
'0' after 80124 ns,
'1' after 80284800 ps,
'0' after 80449600 ps,
'1' after 80692 ns,
'0' after 80774 ns,
'1' after 80855600 ps,
'0' after 80938 ns,
'1' after 81017200 ps,
'0' after 81100400 ps,
'1' after 81180 ns,
'0' after 81264 ns,
'1' after 81342 ns,
'0' after 81425200 ps,
'1' after 81506 ns,
'0' after 81589200 ps,
'1' after 81667600 ps,
'0' after 81750800 ps,
'1' after 81830800 ps,
'0' after 81914400 ps,
'1' after 81993200 ps,
'0' after 82076 ns,
'1' after 82157200 ps,
'0' after 82240 ns,
'1' after 82318 ns,
'0' after 82401600 ps,
'1' after 82482400 ps,
'0' after 82646800 ps,
'1' after 82725600 ps,
'0' after 82809200 ps,
'1' after 82889200 ps,
'0' after 82972800 ps,
'1' after 83132400 ps,
'0' after 83215200 ps,
'1' after 83296400 ps,
'0' after 83378800 ps,
'1' after 83458 ns,
'0' after 83541200 ps,
'1' after 83620800 ps,
'0' after 83704800 ps,
'1' after 83783200 ps,
'0' after 83866400 ps,
'1' after 83947200 ps,
'0' after 84029600 ps,
'1' after 84108800 ps,
'0' after 84192 ns,
'1' after 84272400 ps,
'0' after 84355600 ps,
'1' after 84434 ns,
'0' after 84517200 ps,
'1' after 84598400 ps,
'0' after 84680800 ps,
'1' after 84760400 ps,
'0' after 84843600 ps,
'1' after 84922800 ps,
'0' after 85088400 ps,
'1' after 85166800 ps,
'0' after 85576 ns,
'1' after 85655200 ps,
'0' after 85739600 ps,
'1' after 85816800 ps,
'0' after 85900800 ps,
'1' after 85981200 ps,
'0' after 86064400 ps,
'1' after 86143200 ps,
'0' after 86226400 ps,
'1' after 86306800 ps,
'0' after 86390 ns,
'1' after 86468800 ps,
'0' after 86552 ns,
'1' after 86632 ns,
'0' after 86715600 ps,
'1' after 86794400 ps,
'0' after 86877200 ps,
'1' after 86957600 ps,
'0' after 87041200 ps,
'1' after 87119600 ps,
'0' after 87203200 ps,
'1' after 87283200 ps,
'0' after 87366800 ps,
'1' after 87607600 ps,
'0' after 87772800 ps,
'1' after 88016 ns,
'0' after 88424400 ps,
'1' after 88828 ns,
'0' after 89238 ns,
'1' after 89642800 ps,
'0' after 89970400 ps,
'1' after 90049600 ps,
'0' after 90214400 ps,
'1' after 90292800 ps,
'0' after 90458400 ps,
'1' after 90862400 ps,
'0' after 91272400 ps,
'1' after 91676400 ps,
'0' after 92086 ns,
'1' after 92489600 ps,
'0' after 92573600 ps,
'1' after 92735200 ps,
'0' after 92899200 ps,
'1' after 93304400 ps,
'0' after 93713200 ps,
'1' after 94116800 ps,
'0' after 94527200 ps,
'1' after 94931200 ps,
'0' after 95014 ns,
'1' after 95094400 ps,
'0' after 95178 ns,
'1' after 95256800 ps,
'0' after 95339600 ps,
'1' after 95420400 ps,
'0' after 95503600 ps,
'1' after 95581600 ps,
'0' after 95665200 ps,
'1' after 95745600 ps,
'0' after 95828800 ps,
'1' after 95908 ns,
'0' after 95990400 ps,
'1' after 96070800 ps,
'0' after 96154800 ps,
'1' after 96232400 ps,
'0' after 96316 ns,
'1' after 96396800 ps,
'0' after 96480 ns,
'1' after 96558400 ps,
'0' after 96641200 ps,
'1' after 96722 ns,
'0' after 96805200 ps,
'1' after 96884400 ps,
'0' after 96967200 ps,
'1' after 97047600 ps,
'0' after 97131200 ps,
'1' after 97209600 ps,
'0' after 97374400 ps,
'1' after 97453600 ps,
'0' after 97537600 ps,
'1' after 97616800 ps,
'0' after 97782400 ps,
'1' after 98673200 ps,
'0' after 99084400 ps,
'1' after 99163200 ps,
'0' after 99246400 ps,
'1' after 99326400 ps,
'0' after 99410800 ps,
'1' after 99488800 ps,
'0' after 99571600 ps,
'1' after 99652800 ps,
'0' after 99735600 ps,
'1' after 99814400 ps,
'0' after 99897600 ps,
'1' after 99977600 ps,
'0' after 100061600 ps,
'1' after 100139200 ps,
'0' after 100222400 ps,
'1' after 100304 ns,
'0' after 100386800 ps,
'1' after 100466 ns,
'0' after 100548800 ps,
'1' after 100629200 ps,
'0' after 100712400 ps,
'1' after 100872800 ps,
'0' after 101119600 ps,
'1' after 101523600 ps,
'0' after 101932400 ps,
'1' after 102337600 ps,
'0' after 102746800 ps,
'1' after 103151200 ps,
'0' after 103234 ns,
'1' after 103396400 ps,
'0' after 103560400 ps,
'1' after 103720800 ps,
'0' after 103885600 ps,
'1' after 103965200 ps,
'0' after 104048800 ps,
'1' after 104126800 ps,
'0' after 104210 ns,
'1' after 104291200 ps,
'0' after 104373600 ps,
'1' after 104452800 ps,
'0' after 104535600 ps,
'1' after 104616400 ps,
'0' after 104699600 ps,
'1' after 104778400 ps,
'0' after 104861200 ps,
'1' after 104942400 ps,
'0' after 105024800 ps,
'1' after 105103600 ps,
'0' after 105187200 ps,
'1' after 105267200 ps,
'0' after 105351200 ps,
'1' after 105428400 ps,
'0' after 105511600 ps,
'1' after 105593200 ps,
'0' after 105676 ns,
'1' after 105754800 ps,
'0' after 105838 ns,
'1' after 105918 ns,
'0' after 106002 ns,
'1' after 106079600 ps,
'0' after 106245200 ps,
'1' after 106406800 ps,
'0' after 106489600 ps,
'1' after 106568 ns,
'0' after 106651600 ps,
'1' after 106732 ns,
'0' after 106815200 ps,
'1' after 106893600 ps,
'0' after 106977200 ps,
'1' after 107058 ns,
'0' after 107140400 ps,
'1' after 107219200 ps,
'0' after 107302400 ps,
'1' after 107383200 ps,
'0' after 107466 ns,
'1' after 107544800 ps,
'0' after 107627600 ps,
'1' after 107708800 ps,
'0' after 107791600 ps,
'1' after 107870800 ps,
'0' after 107953600 ps,
'1' after 108034 ns,
'0' after 108117200 ps,
'1' after 108277200 ps,
'0' after 108360 ns,
'1' after 108440800 ps,
'0' after 108605600 ps,
'1' after 108684 ns,
'0' after 108849200 ps,
'1' after 108928400 ps,
'0' after 109012 ns,
'1' after 109091200 ps,
'0' after 109174800 ps,
'1' after 109254 ns,
'0' after 109338 ns,
'1' after 109415200 ps,
'0' after 109499600 ps,
'1' after 109580 ns,
'0' after 109663200 ps,
'1' after 109741600 ps,
'0' after 109825200 ps,
'1' after 109905600 ps,
'0' after 109988800 ps,
'1' after 110067600 ps,
'0' after 110150800 ps,
'1' after 110231200 ps,
'0' after 110314400 ps,
'1' after 110392 ns,
'0' after 110476 ns,
'1' after 110556800 ps,
'0' after 110802400 ps,
'1' after 110882 ns,
'0' after 111046400 ps,
'1' after 111125200 ps,
'0' after 111208400 ps,
'1' after 111288800 ps,
'0' after 111372400 ps,
'1' after 111450400 ps,
'0' after 111533600 ps,
'1' after 111614 ns,
'0' after 111697200 ps,
'1' after 111776400 ps,
'0' after 111859200 ps,
'1' after 111939600 ps,
'0' after 112022800 ps,
'1' after 112101600 ps,
'0' after 112184400 ps,
'1' after 112265200 ps,
'0' after 112348 ns,
'1' after 112427200 ps,
'0' after 112510800 ps,
'1' after 112590 ns,
'0' after 112674400 ps,
'1' after 112752400 ps,
'0' after 112835600 ps,
'1' after 112916400 ps,
'0' after 112999200 ps,
'1' after 113078 ns,
'0' after 113243200 ps,
'1' after 113322400 ps,
'0' after 113487600 ps,
'1' after 113566 ns,
'0' after 113649600 ps,
'1' after 113729600 ps,
'0' after 114138800 ps,
'1' after 114542800 ps,
'0' after 114952400 ps,
'1' after 115356 ns,
'0' after 115684400 ps,
'1' after 115763200 ps,
'0' after 115846400 ps,
'1' after 115926800 ps,
'0' after 116091200 ps,
'1' after 116170 ns,
'0' after 116170400 ps,
'1' after 116170800 ps,
'0' after 116579600 ps,
'1' after 116984 ns,
'0' after 117393600 ps,
'1' after 117797600 ps,
'0' after 118125600 ps,
'1' after 118204400 ps,
'0' after 118370 ns,
'1' after 118530 ns,
'0' after 118612800 ps,
'1' after 119506400 ps,
'0' after 119916400 ps,
'1' after 119995600 ps,
'0' after 120078800 ps,
'1' after 120158400 ps,
'0' after 120242400 ps,
'1' after 120320800 ps,
'0' after 120404 ns,
'1' after 120484 ns,
'0' after 120568 ns,
'1' after 120646 ns,
'0' after 120729200 ps,
'1' after 120810 ns,
'0' after 120893200 ps,
'1' after 120972 ns,
'0' after 121055200 ps,
'1' after 121135600 ps,
'0' after 121219200 ps,
'1' after 121298 ns,
'0' after 121380400 ps,
'1' after 121461200 ps,
'0' after 121544400 ps,
'1' after 121705200 ps,
'0' after 121788 ns,
'1' after 121950 ns,
'0' after 122357600 ps,
'1' after 122436800 ps,
'0' after 122521200 ps,
'1' after 122599200 ps,
'0' after 122682800 ps,
'1' after 122763200 ps,
'0' after 122846800 ps,
'1' after 122924800 ps,
'0' after 123008 ns,
'1' after 123088800 ps,
'0' after 123172 ns,
'1' after 123250800 ps,
'0' after 123334 ns,
'1' after 123413600 ps,
'0' after 123498 ns,
'1' after 123575600 ps,
'0' after 123658800 ps,
'1' after 123740400 ps,
'0' after 123822800 ps,
'1' after 123902 ns,
'0' after 123985600 ps,
'1' after 124064400 ps,
'0' after 124230 ns,
'1' after 124390400 ps,
'0' after 124473200 ps,
'1' after 124553200 ps,
'0' after 124636800 ps,
'1' after 124714800 ps,
'0' after 124798400 ps,
'1' after 125204400 ps,
'0' after 125613200 ps,
'1' after 126017600 ps,
'0' after 126426800 ps,
'1' after 126587200 ps,
'0' after 126752 ns,
'1' after 126831200 ps,
'0' after 126914800 ps,
'1' after 126992800 ps,
'0' after 127240400 ps,
'1' after 127318800 ps,
'0' after 127402400 ps,
'1' after 127482 ns,
'0' after 127566400 ps,
'1' after 127644 ns,
'0' after 127727600 ps,
'1' after 127808400 ps,
'0' after 127891200 ps,
'1' after 127969600 ps,
'0' after 128053600 ps,
'1' after 128134 ns,
'0' after 128217200 ps,
'1' after 128294800 ps,
'0' after 128378400 ps,
'1' after 128459600 ps,
'0' after 128542400 ps,
'1' after 128620800 ps,
'0' after 128704 ns,
'1' after 128784800 ps,
'0' after 128868 ns,
'1' after 128946 ns,
'0' after 128946400 ps,
'1' after 128946800 ps,
'0' after 129030 ns,
'1' after 129110 ns,
'0' after 129193600 ps,
'1' after 129271200 ps,
'0' after 129354800 ps,
'1' after 129517600 ps,
'0' after 129681200 ps,
'1' after 130086400 ps,
'0' after 130495200 ps,
'1' after 130898800 ps,
'0' after 131309200 ps,
'1' after 131631600 ps,
'0' after 131714 ns,
'1' after 131795600 ps,
'0' after 132122800 ps,
'1' after 132526400 ps,
'0' after 132936400 ps,
'1' after 133340400 ps,
'0' after 133749600 ps,
'1' after 133992 ns,
'0' after 134074400 ps,
'1' after 134155600 ps,
'0' after 134400800 ps,
'1' after 134561600 ps,
'0' after 134970800 ps,
'1' after 135374800 ps,
'0' after 135784 ns,
'1' after 136188400 ps,
'0' after 136435200 ps,
'1' after 136514400 ps,
'0' after 136597200 ps,
'1' after 136759200 ps,
'0' after 137004800 ps,
'1' after 137083600 ps,
'0' after 137168 ns,
'1' after 137246 ns,
'0' after 137329200 ps,
'1' after 137409600 ps,
'0' after 137493200 ps,
'1' after 137571200 ps,
'0' after 137654800 ps,
'1' after 137735600 ps,
'0' after 137818400 ps,
'1' after 137897200 ps,
'0' after 137980400 ps,
'1' after 138060800 ps,
'0' after 138144400 ps,
'1' after 138222800 ps,
'0' after 138305600 ps,
'1' after 138386400 ps,
'0' after 138470 ns,
'1' after 138548400 ps,
'0' after 138631200 ps,
'1' after 138712 ns,
'0' after 138795200 ps,
'1' after 138873200 ps,
'0' after 139038800 ps,
'1' after 139444 ns,
'0' after 140341200 ps,
'1' after 140745600 ps,
'0' after 140829200 ps,
'1' after 140909200 ps,
'0' after 140992400 ps,
'1' after 141072 ns,
'0' after 141154800 ps,
'1' after 141235600 ps,
'0' after 141318400 ps,
'1' after 141397600 ps,
'0' after 141480400 ps,
'1' after 141561200 ps,
'0' after 141644 ns,
'1' after 141722800 ps,
'0' after 141806 ns,
'1' after 141886800 ps,
'0' after 141969600 ps,
'1' after 142048400 ps,
'0' after 142131200 ps,
'1' after 142212400 ps,
'0' after 142295200 ps,
'1' after 142373600 ps,
'0' after 142456800 ps,
'1' after 142537600 ps,
'0' after 142620400 ps,
'1' after 142781200 ps,
'0' after 142945200 ps,
'1' after 143188800 ps,
'0' after 143597200 ps,
'1' after 144001200 ps,
'0' after 144410800 ps,
'1' after 144814800 ps,
'0' after 145224800 ps,
'1' after 145467200 ps,
'0' after 145549200 ps,
'1' after 145630 ns,
'0' after 145712800 ps,
'1' after 145791600 ps,
'0' after 145874800 ps,
'1' after 145954800 ps,
'0' after 145955200 ps,
'1' after 145955600 ps,
'0' after 146038400 ps,
'1' after 146117200 ps,
'0' after 146199600 ps,
'1' after 146280800 ps,
'0' after 146364 ns,
'1' after 146442400 ps,
'0' after 146525600 ps,
'1' after 146606 ns,
'0' after 146689600 ps,
'1' after 146767600 ps,
'0' after 146850800 ps,
'1' after 146931200 ps,
'0' after 147014800 ps,
'1' after 147093200 ps,
'0' after 147176400 ps,
'1' after 147257200 ps,
'0' after 147340 ns,
'1' after 147419600 ps,
'0' after 147665600 ps,
'1' after 147744 ns,
'0' after 148072800 ps,
'1' after 148476400 ps,
'0' after 148886400 ps,
'1' after 149290400 ps,
'0' after 149700 ns,
'1' after 150103600 ps,
'0' after 150513600 ps,
'1' after 150918 ns,
'0' after 151327200 ps,
'1' after 151731200 ps,
'0' after 152140800 ps,
'1' after 152301600 ps,
'0' after 152548 ns,
'1' after 152789600 ps,
'0' after 152872 ns,
'1' after 152953200 ps,
'0' after 153035600 ps,
'1' after 153114800 ps,
'0' after 153198400 ps,
'1' after 153278 ns,
'0' after 153362 ns,
'1' after 153440 ns,
'0' after 153523200 ps,
'1' after 153604 ns,
'0' after 153686800 ps,
'1' after 153766 ns,
'0' after 153849200 ps,
'1' after 153929600 ps,
'0' after 154012800 ps,
'1' after 154090400 ps,
'0' after 154174400 ps,
'1' after 154254400 ps,
'0' after 154338 ns,
'1' after 154416800 ps,
'0' after 154499600 ps,
'1' after 154580 ns,
'0' after 154663600 ps,
'1' after 154742 ns,
'0' after 154824800 ps,
'1' after 154906 ns,
'0' after 154988800 ps,
'1' after 155067200 ps,
'0' after 155314800 ps,
'1' after 155393200 ps,
'0' after 155476800 ps,
'1' after 155556800 ps,
'0' after 155640 ns,
'1' after 155718400 ps,
'0' after 155801600 ps,
'1' after 155882 ns,
'0' after 155965600 ps,
'1' after 156044 ns,
'0' after 156127200 ps,
'1' after 156208 ns,
'0' after 156290800 ps,
'1' after 156369600 ps,
'0' after 156452800 ps,
'1' after 156532800 ps,
'0' after 156616800 ps,
'1' after 156695200 ps,
'0' after 156778400 ps,
'1' after 156858800 ps,
'0' after 156942 ns,
'1' after 157020400 ps,
'0' after 157103600 ps,
'1' after 157265200 ps,
'0' after 157349200 ps,
'1' after 157427200 ps,
'0' after 157837200 ps,
'1' after 158241200 ps,
'0' after 158650800 ps,
'1' after 159056 ns,
'0' after 159464800 ps,
'1' after 159868400 ps,
'0' after 160034 ns,
'1' after 160276 ns,
'0' after 161173600 ps,
'1' after 161578 ns,
'0' after 161988 ns,
'1' after 162392 ns,
'0' after 162801600 ps,
'1' after 163205600 ps,
'0' after 163289200 ps,
'1' after 163369600 ps,
'0' after 163615600 ps,
'1' after 164019600 ps,
'0' after 164102 ns,
'1' after 164183600 ps,
'0' after 164266400 ps,
'1' after 164345200 ps,
'0' after 164428 ns,
'1' after 164508800 ps,
'0' after 164592400 ps,
'1' after 164670400 ps,
'0' after 164753600 ps,
'1' after 164834800 ps,
'0' after 164917200 ps,
'1' after 164996 ns,
'0' after 165079200 ps,
'1' after 165159600 ps,
'0' after 165242800 ps,
'1' after 165321200 ps,
'0' after 165404 ns,
'1' after 165486 ns,
'0' after 165568 ns,
'1' after 165647600 ps,
'0' after 165730800 ps,
'1' after 165810400 ps,
'0' after 166056400 ps,
'1' after 166135600 ps,
'0' after 166382400 ps,
'1' after 166460800 ps,
'0' after 166543600 ps,
'1' after 166624 ns,
'0' after 166708 ns,
'1' after 166785600 ps,
'0' after 166869200 ps,
'1' after 166950 ns,
'0' after 167032800 ps,
'1' after 167111600 ps,
'0' after 167195200 ps,
'1' after 167275200 ps,
'0' after 167358800 ps,
'1' after 167437200 ps,
'0' after 167520400 ps,
'1' after 167600800 ps,
'0' after 167684 ns,
'1' after 167762800 ps,
'0' after 167846 ns,
'1' after 167926400 ps,
'0' after 168009600 ps,
'1' after 168088400 ps,
'0' after 168171200 ps,
'1' after 168252 ns,
'0' after 168416400 ps,
'1' after 168494800 ps,
'0' after 168904400 ps,
'1' after 168983200 ps,
'0' after 169066800 ps,
'1' after 169146400 ps,
'0' after 169230400 ps,
'1' after 169308400 ps,
'0' after 169391600 ps,
'1' after 169472800 ps,
'0' after 169555200 ps,
'1' after 169634400 ps,
'0' after 169719200 ps,
'1' after 169796800 ps,
'0' after 169879600 ps,
'1' after 169961200 ps,
'0' after 170043600 ps,
'1' after 170122800 ps,
'0' after 170206800 ps,
'1' after 170285200 ps,
'0' after 170368400 ps,
'1' after 170448800 ps,
'0' after 170532 ns,
'1' after 170610800 ps,
'0' after 170693600 ps,
'1' after 170937200 ps,
'0' after 171264400 ps,
'1' after 171342800 ps,
'0' after 171752800 ps,
'1' after 172156800 ps,
'0' after 172566 ns,
'1' after 172970800 ps,
'0' after 173299200 ps,
'1' after 173377200 ps,
'0' after 173461200 ps,
'1' after 173539600 ps,
'0' after 173705200 ps,
'1' after 173784 ns,
'0' after 174193200 ps,
'1' after 174598400 ps,
'0' after 175007600 ps,
'1' after 175412 ns,
'0' after 175820400 ps,
'1' after 175900400 ps,
'0' after 176065200 ps,
'1' after 176143600 ps,
'0' after 176227600 ps,
'1' after 176632400 ps,
'0' after 177042400 ps,
'1' after 177445600 ps,
'0' after 177855600 ps,
'1' after 178016 ns,
'0' after 178262 ns,
'1' after 178422800 ps,
'0' after 178505200 ps,
'1' after 178586 ns,
'0' after 178669200 ps,
'1' after 178747600 ps,
'0' after 178830800 ps,
'1' after 178911600 ps,
'0' after 178994800 ps,
'1' after 179072800 ps,
'0' after 179156800 ps,
'1' after 179236800 ps,
'0' after 179320400 ps,
'1' after 179398800 ps,
'0' after 179482 ns,
'1' after 179562800 ps,
'0' after 179645600 ps,
'1' after 179724 ns,
'0' after 179807600 ps,
'1' after 179887600 ps,
'0' after 179971200 ps,
'1' after 180049600 ps,
'0' after 180132800 ps,
'1' after 180213200 ps,
'0' after 180296400 ps,
'1' after 180375200 ps,
'0' after 180458400 ps,
'1' after 180538800 ps,
'0' after 180622 ns,
'1' after 180700800 ps,
'0' after 180784 ns,
'1' after 180864400 ps,
'0' after 181028800 ps,
'1' after 181108400 ps,
'0' after 182006 ns,
'1' after 182410 ns,
'0' after 182493200 ps,
'1' after 182574400 ps,
'0' after 182657200 ps,
'1' after 182736 ns,
'0' after 182820400 ps,
'1' after 182898400 ps,
'0' after 182982 ns,
'1' after 183062400 ps,
'0' after 183146 ns,
'1' after 183224400 ps,
'0' after 183307200 ps,
'1' after 183388400 ps,
'0' after 183471200 ps,
'1' after 183549600 ps,
'0' after 183632800 ps,
'1' after 183713600 ps,
'0' after 183796800 ps,
'1' after 183874800 ps,
'0' after 183958 ns,
'1' after 184039600 ps,
'0' after 184122400 ps,
'1' after 184200800 ps,
'0' after 184366 ns,
'1' after 184445200 ps,
'0' after 184610 ns,
'1' after 184689200 ps,
'0' after 184854400 ps,
'1' after 184933600 ps,
'0' after 185016800 ps,
'1' after 185096 ns,
'0' after 185180400 ps,
'1' after 185258400 ps,
'0' after 185341600 ps,
'1' after 185422400 ps,
'0' after 185505600 ps,
'1' after 185584400 ps,
'0' after 185667600 ps,
'1' after 185748 ns,
'0' after 185831200 ps,
'1' after 185909200 ps,
'0' after 185992800 ps,
'1' after 186073200 ps,
'0' after 186156400 ps,
'1' after 186234400 ps,
'0' after 186318 ns,
'1' after 186399200 ps,
'0' after 186481600 ps,
'1' after 186642400 ps,
'0' after 186724800 ps,
'1' after 186806 ns,
'0' after 186888800 ps,
'1' after 187049200 ps,
'0' after 187296 ns,
'1' after 187700400 ps,
'0' after 188109600 ps,
'1' after 188513200 ps,
'0' after 188923200 ps,
'1' after 189164800 ps,
'0' after 189247200 ps,
'1' after 189328400 ps,
'0' after 189410800 ps,
'1' after 189571600 ps,
'0' after 189654 ns,
'1' after 189735200 ps,
'0' after 189818 ns,
'1' after 189897200 ps,
'0' after 189980 ns,
'1' after 190060400 ps,
'0' after 190143600 ps,
'1' after 190222 ns,
'0' after 190304800 ps,
'1' after 190386 ns,
'0' after 190468800 ps,
'1' after 190548 ns,
'0' after 190631200 ps,
'1' after 190710800 ps,
'0' after 190794400 ps,
'1' after 190873200 ps,
'0' after 190956 ns,
'1' after 191036800 ps,
'0' after 191120 ns,
'1' after 191198800 ps,
'0' after 191281600 ps,
'1' after 191362800 ps,
'0' after 191445200 ps,
'1' after 191768400 ps,
'0' after 191851200 ps,
'1' after 192014 ns,
'0' after 192177600 ps,
'1' after 192582400 ps,
'0' after 192991200 ps,
'1' after 193395600 ps,
'0' after 193805200 ps,
'1' after 194128400 ps,
'0' after 194210400 ps,
'1' after 194373600 ps,
'0' after 194456400 ps,
'1' after 194616400 ps,
'0' after 194698800 ps,
'1' after 194780800 ps,
'0' after 194862800 ps,
'1' after 194942400 ps,
'0' after 195025200 ps,
'1' after 195104800 ps,
'0' after 195188 ns,
'1' after 195267600 ps,
'0' after 195351200 ps,
'1' after 195430 ns,
'0' after 195512800 ps,
'1' after 195594 ns,
'0' after 195676800 ps,
'1' after 195756 ns,
'0' after 195838800 ps,
'1' after 195918800 ps,
'0' after 196002400 ps,
'1' after 196080800 ps,
'0' after 196163600 ps,
'1' after 196244800 ps,
'0' after 196327200 ps,
'1' after 196406400 ps,
'0' after 196490 ns,
'1' after 196651200 ps,
'0' after 196733600 ps,
'1' after 196814 ns,
'0' after 197060 ns,
'1' after 197464800 ps,
'0' after 197873600 ps,
'1' after 198278 ns,
'0' after 198687600 ps,
'1' after 199010800 ps,
'0' after 199093200 ps,
'1' after 199418800 ps,
'0' after 199500 ns,
'1' after 199906 ns,
'0' after 200314800 ps,
'1' after 200718800 ps,
'0' after 201128400 ps,
'1' after 201370400 ps,
'0' after 201534400 ps,
'1' after 201696800 ps,
'0' after 201942 ns,
'1' after 202834 ns,
'0' after 203245200 ps,
'1' after 203324400 ps,
'0' after 203406800 ps,
'1' after 203486800 ps,
'0' after 203570400 ps,
'1' after 203649200 ps,
'0' after 203732400 ps,
'1' after 203812800 ps,
'0' after 203896400 ps,
'1' after 203974400 ps,
'0' after 204057600 ps,
'1' after 204138400 ps,
'0' after 204221600 ps,
'1' after 204300400 ps,
'0' after 204383200 ps,
'1' after 204463600 ps,
'0' after 204547200 ps,
'1' after 204626 ns,
'0' after 204708800 ps,
'1' after 204789200 ps,
'0' after 204872800 ps,
'1' after 204951600 ps,
'0' after 205034800 ps,
'1' after 205278 ns,
'0' after 205359600 ps,
'1' after 205604 ns,
'0' after 205684800 ps,
'1' after 205766 ns,
'0' after 205849600 ps,
'1' after 205928 ns,
'0' after 206010800 ps,
'1' after 206091200 ps,
'0' after 206174800 ps,
'1' after 206253200 ps,
'0' after 206336400 ps,
'1' after 206416800 ps,
'0' after 206500400 ps,
'1' after 206578800 ps,
'0' after 206662 ns,
'1' after 206742800 ps,
'0' after 206825600 ps,
'1' after 206904 ns,
'0' after 206987200 ps,
'1' after 207068 ns,
'0' after 207150800 ps,
'1' after 207229600 ps,
'0' after 207312800 ps,
'1' after 207393600 ps,
'0' after 207476800 ps,
'1' after 207718 ns,
'0' after 207801200 ps,
'1' after 208126400 ps,
'0' after 208534400 ps,
'1' after 208938800 ps,
'0' after 209347600 ps,
'1' after 209752400 ps,
'0' after 210080400 ps,
'1' after 210158800 ps,
'0' after 210242800 ps,
'1' after 210566400 ps,
'0' after 210648400 ps,
'1' after 210730400 ps,
'0' after 210812400 ps,
'1' after 210891200 ps,
'0' after 210974400 ps,
'1' after 211054400 ps,
'0' after 211138400 ps,
'1' after 211216400 ps,
'0' after 211299600 ps,
'1' after 211381200 ps,
'0' after 211463200 ps,
'1' after 211542400 ps,
'0' after 211625600 ps,
'1' after 211706400 ps,
'0' after 211790 ns,
'1' after 211867200 ps,
'0' after 211950400 ps,
'1' after 212031600 ps,
'0' after 212114800 ps,
'1' after 212193600 ps,
'0' after 212276400 ps,
'1' after 212356800 ps,
'0' after 212602800 ps,
'1' after 212682 ns,
'0' after 212766 ns,
'1' after 213007600 ps,
'0' after 213090 ns,
'1' after 213171200 ps,
'0' after 213253600 ps,
'1' after 213332400 ps,
'0' after 213415600 ps,
'1' after 213496400 ps,
'0' after 213579200 ps,
'1' after 213657600 ps,
'0' after 213740800 ps,
'1' after 213822 ns,
'0' after 213904800 ps,
'1' after 213983600 ps,
'0' after 214066800 ps,
'1' after 214146800 ps,
'0' after 214230 ns,
'1' after 214308800 ps,
'0' after 214392 ns,
'1' after 214472800 ps,
'0' after 214556 ns,
'1' after 214634800 ps,
'0' after 214717200 ps,
'1' after 214798400 ps,
'0' after 214881200 ps,
'1' after 214960 ns,
'0' after 215043600 ps,
'1' after 215205200 ps,
'0' after 215287600 ps,
'1' after 215449200 ps,
'0' after 215857600 ps,
'1' after 216262 ns,
'0' after 216670800 ps,
'1' after 217075600 ps,
'0' after 217240400 ps,
'1' after 217320400 ps,
'0' after 217404 ns,
'1' after 217481600 ps,
'0' after 217565600 ps,
'1' after 217890 ns,
'0' after 217890400 ps,
'1' after 217890800 ps,
'0' after 217972 ns,
'1' after 218053200 ps,
'0' after 218135600 ps,
'1' after 218214800 ps,
'0' after 218298400 ps,
'1' after 218378 ns,
'0' after 218462 ns,
'1' after 218540 ns,
'0' after 218623200 ps,
'1' after 218703600 ps,
'0' after 218704 ns,
'1' after 218704400 ps,
'0' after 218787200 ps,
'1' after 218866400 ps,
'0' after 218949200 ps,
'1' after 219029200 ps,
'0' after 219112400 ps,
'1' after 219191200 ps,
'0' after 219274400 ps,
'1' after 219355200 ps,
'0' after 219437600 ps,
'1' after 219517200 ps,
'0' after 219600 ns,
'1' after 219680 ns,
'0' after 219926400 ps,
'1' after 220005200 ps,
'0' after 220088400 ps,
'1' after 220331200 ps,
'0' after 220740 ns,
'1' after 221144 ns,
'0' after 221554 ns,
'1' after 221958 ns,
'0' after 222367600 ps,
'1' after 222690400 ps,
'0' after 222773600 ps,
'1' after 223666800 ps,
'0' after 224077200 ps,
'1' after 224481200 ps,
'0' after 224890800 ps,
'1' after 225295200 ps,
'0' after 225704800 ps,
'1' after 226109200 ps,
'0' after 226192 ns,
'1' after 226354 ns,
'0' after 226436 ns,
'1' after 226516400 ps,
'0' after 226925200 ps,
'1' after 227330 ns,
'0' after 227739200 ps,
'1' after 228143200 ps,
'0' after 228390 ns,
'1' after 228469600 ps,
'0' after 228552400 ps,
'1' after 228631600 ps,
'0' after 228714400 ps,
'1' after 228795200 ps,
'0' after 228878400 ps,
'1' after 228957200 ps,
'0' after 229040400 ps,
'1' after 229120800 ps,
'0' after 229203600 ps,
'1' after 229282400 ps,
'0' after 229365600 ps,
'1' after 229446400 ps,
'0' after 229529200 ps,
'1' after 229607600 ps,
'0' after 229690800 ps,
'1' after 229771600 ps,
'0' after 229854800 ps,
'1' after 229933600 ps,
'0' after 230016400 ps,
'1' after 230097600 ps,
'0' after 230180400 ps,
'1' after 230259200 ps,
'0' after 230342400 ps,
'1' after 230422400 ps,
'0' after 230505600 ps,
'1' after 230584 ns,
'0' after 230667600 ps,
'1' after 230748400 ps,
'0' after 230912400 ps,
'1' after 230992 ns,
'0' after 231075200 ps,
'1' after 231235600 ps,
'0' after 231400400 ps,
'1' after 231805200 ps,
'0' after 232214800 ps,
'1' after 232618800 ps,
'0' after 233028 ns,
'1' after 233351200 ps,
'0' after 233433200 ps,
'1' after 233597200 ps,
'0' after 233679200 ps,
'1' after 233839600 ps,
'0' after 234248800 ps,
'1' after 234652800 ps,
'0' after 235062400 ps,
'1' after 235466400 ps,
'0' after 235631600 ps,
'1' after 235792800 ps,
'0' after 235875200 ps,
'1' after 235955600 ps,
'0' after 236120 ns,
'1' after 236199600 ps,
'0' after 236282800 ps,
'1' after 236687200 ps,
'0' after 237096400 ps,
'1' after 237501200 ps,
'0' after 237910400 ps,
'1' after 238071200 ps,
'0' after 238235600 ps,
'1' after 238314800 ps,
'0' after 238724400 ps,
'1' after 238802800 ps,
'0' after 238886 ns,
'1' after 238966 ns,
'0' after 239050 ns,
'1' after 239127600 ps,
'0' after 239211200 ps,
'1' after 239292400 ps,
'0' after 239375200 ps,
'1' after 239453600 ps,
'0' after 239537200 ps,
'1' after 239617200 ps,
'0' after 239701200 ps,
'1' after 239779200 ps,
'0' after 239862 ns,
'1' after 239942800 ps,
'0' after 240026400 ps,
'1' after 240104800 ps,
'0' after 240188 ns,
'1' after 240268400 ps,
'0' after 240352 ns,
'1' after 240430 ns,
'0' after 240513200 ps,
'1' after 240594 ns,
'0' after 240677200 ps,
'1' after 240756 ns,
'0' after 240838800 ps,
'1' after 241001200 ps,
'0' after 241164800 ps,
'1' after 241569200 ps,
'0' after 241978800 ps,
'1' after 242383200 ps,
'0' after 242793200 ps,
'1' after 243115600 ps,
'0' after 243198 ns,
'1' after 243278800 ps,
'0' after 243362 ns,
'1' after 243440400 ps,
'0' after 243524400 ps,
'1' after 243604800 ps,
'0' after 244501600 ps,
'1' after 244906400 ps,
'0' after 244989600 ps,
'1' after 245070 ns,
'0' after 245153200 ps,
'1' after 245232 ns,
'0' after 245315200 ps,
'1' after 245395600 ps,
'0' after 245478800 ps,
'1' after 245557600 ps,
'0' after 245640800 ps,
'1' after 245721200 ps,
'0' after 245804800 ps,
'1' after 245883200 ps,
'0' after 245966 ns,
'1' after 246047200 ps,
'0' after 246130 ns,
'1' after 246208400 ps,
'0' after 246291600 ps,
'1' after 246372400 ps,
'0' after 246455600 ps,
'1' after 246534 ns,
'0' after 246617200 ps,
'1' after 246697600 ps,
'0' after 246943600 ps,
'1' after 247022800 ps,
'0' after 247106800 ps,
'1' after 247184800 ps,
'0' after 247268 ns,
'1' after 247349200 ps,
'0' after 247757600 ps,
'1' after 248162 ns,
'0' after 248571600 ps,
'1' after 248975200 ps,
'0' after 249222400 ps,
'1' after 249300800 ps,
'0' after 249384800 ps,
'1' after 249708400 ps,
'0' after 249790800 ps,
'1' after 249871600 ps,
'0' after 249954400 ps,
'1' after 250033600 ps,
'0' after 250116400 ps,
'1' after 250196800 ps,
'0' after 250280400 ps,
'1' after 250359200 ps,
'0' after 250441600 ps,
'1' after 250522400 ps,
'0' after 250605200 ps,
'1' after 250684 ns,
'0' after 250767600 ps,
'1' after 250847600 ps,
'0' after 250931200 ps,
'1' after 251009200 ps,
'0' after 251092400 ps,
'1' after 251174 ns,
'0' after 251256400 ps,
'1' after 251335200 ps,
'0' after 251418 ns,
'1' after 251580 ns,
'0' after 251663200 ps,
'1' after 251823600 ps,
'0' after 251906 ns,
'1' after 251987200 ps,
'0' after 252070 ns,
'1' after 252230800 ps,
'0' after 252639600 ps,
'1' after 253044400 ps,
'0' after 253453200 ps,
'1' after 253858 ns,
'0' after 254266800 ps,
'1' after 254346 ns,
'0' after 254674 ns,
'1' after 254752800 ps,
'0' after 254836 ns,
'1' after 254915600 ps,
'0' after 255 us,
'1' after 255077600 ps,
'0' after 255160800 ps,
'1' after 255242 ns,
'0' after 255324800 ps,
'1' after 255403600 ps,
'0' after 255487200 ps,
'1' after 255566400 ps,
'0' after 255651200 ps,
'1' after 255728800 ps,
'0' after 255812 ns,
'1' after 255892800 ps,
'0' after 255976 ns,
'1' after 256054800 ps,
'0' after 256137600 ps,
'1' after 256218400 ps,
'0' after 256301600 ps,
'1' after 256461600 ps,
'0' after 256544400 ps,
'1' after 256625200 ps,
'0' after 256708400 ps,
'1' after 256786800 ps,
'0' after 256870 ns,
'1' after 257113600 ps,
'0' after 257195200 ps,
'1' after 257275600 ps,
'0' after 257359200 ps,
'1' after 257437600 ps,
'0' after 257520800 ps,
'1' after 257602 ns,
'0' after 257684400 ps,
'1' after 257763600 ps,
'0' after 257846800 ps,
'1' after 257927200 ps,
'0' after 258010800 ps,
'1' after 258088400 ps,
'0' after 258171200 ps,
'1' after 258253200 ps,
'0' after 258335600 ps,
'1' after 258414400 ps,
'0' after 258497200 ps,
'1' after 258578400 ps,
'0' after 258661200 ps,
'1' after 258740 ns,
'0' after 258822400 ps,
'1' after 259147600 ps,
'0' after 259229600 ps,
'1' after 259392 ns,
'0' after 259556400 ps,
'1' after 259960400 ps,
'0' after 260370 ns,
'1' after 260773600 ps,
'0' after 261183600 ps,
'1' after 261587600 ps,
'0' after 261670400 ps,
'1' after 261751600 ps,
'0' after 261834 ns,
'1' after 261914 ns,
'0' after 261997200 ps,
'1' after 262076400 ps,
'0' after 262159600 ps,
'1' after 262239600 ps,
'0' after 262323200 ps,
'1' after 262400800 ps,
'0' after 262484800 ps,
'1' after 262566 ns,
'0' after 262648 ns,
'1' after 262727200 ps,
'0' after 262810400 ps,
'1' after 262890400 ps,
'0' after 262974 ns,
'1' after 263052 ns,
'0' after 263135200 ps,
'1' after 263216400 ps,
'0' after 263298400 ps,
'1' after 263378400 ps,
'0' after 263462800 ps,
'1' after 263540400 ps,
'0' after 263623600 ps,
'1' after 263704800 ps,
'0' after 263787200 ps,
'1' after 263866 ns,
'0' after 264031200 ps,
'1' after 264110400 ps,
'0' after 264194400 ps,
'1' after 264274 ns,
'0' after 264438400 ps,
'1' after 265329600 ps,
'0' after 265741200 ps,
'1' after 266145600 ps,
'0' after 266554800 ps,
'1' after 266959200 ps,
'0' after 267369200 ps,
'1' after 267692800 ps,
'0' after 267774400 ps,
'1' after 268100 ns,
'0' after 268181600 ps,
'1' after 268262400 ps,
'0' after 268345600 ps,
'1' after 268424400 ps,
'0' after 268506800 ps,
'1' after 268588 ns,
'0' after 268670800 ps,
'1' after 268750 ns,
'0' after 268832400 ps,
'1' after 268912800 ps,
'0' after 268996800 ps,
'1' after 269075200 ps,
'0' after 269158 ns,
'1' after 269238800 ps,
'0' after 269322 ns,
'1' after 269400800 ps,
'0' after 269483200 ps,
'1' after 269564400 ps,
'0' after 269647600 ps,
'1' after 269726400 ps,
'0' after 269809200 ps,
'1' after 269889600 ps,
'0' after 270054800 ps,
'1' after 270214800 ps,
'0' after 270296800 ps,
'1' after 270378800 ps,
'0' after 270542400 ps,
'1' after 270621600 ps,
'0' after 271030800 ps,
'1' after 271434400 ps,
'0' after 271844400 ps,
'1' after 272248800 ps,
'0' after 272495200 ps,
'1' after 272656 ns,
'0' after 272820400 ps,
'1' after 272900 ns,
'0' after 273064800 ps,
'1' after 273144 ns,
'0' after 273227200 ps,
'1' after 273306400 ps,
'0' after 273390400 ps,
'1' after 273468800 ps,
'0' after 273552400 ps,
'1' after 273632400 ps,
'0' after 273716400 ps,
'1' after 273794400 ps,
'0' after 273878 ns,
'1' after 273958400 ps,
'0' after 274041600 ps,
'1' after 274119600 ps,
'0' after 274203200 ps,
'1' after 274284 ns,
'0' after 274366800 ps,
'1' after 274446 ns,
'0' after 274528800 ps,
'1' after 274609600 ps,
'0' after 274692 ns,
'1' after 274771200 ps,
'0' after 274936 ns,
'1' after 275097200 ps,
'0' after 275179600 ps,
'1' after 275504400 ps,
'0' after 275913200 ps,
'1' after 276317200 ps,
'0' after 276726400 ps,
'1' after 277131200 ps,
'0' after 277540 ns,
'1' after 277700800 ps,
'0' after 277947200 ps,
'1' after 278025600 ps,
'0' after 278109200 ps,
'1' after 278189200 ps,
'0' after 278273200 ps,
'1' after 278351200 ps,
'0' after 278434400 ps,
'1' after 278515200 ps,
'0' after 278598 ns,
'1' after 278676800 ps,
'0' after 278760400 ps,
'1' after 278840400 ps,
'0' after 278924 ns,
'1' after 279002 ns,
'0' after 279085200 ps,
'1' after 279166800 ps,
'0' after 279248800 ps,
'1' after 279328 ns,
'0' after 279411600 ps,
'1' after 279490800 ps,
'0' after 279575200 ps,
'1' after 279652800 ps,
'0' after 279981600 ps,
'1' after 280060400 ps,
'0' after 280225200 ps,
'1' after 280386400 ps,
'0' after 280795600 ps,
'1' after 281199600 ps,
'0' after 281608800 ps,
'1' after 282013200 ps,
'0' after 282341600 ps,
'1' after 282420 ns,
'0' after 282504 ns,
'1' after 282827600 ps,
'0' after 282909200 ps,
'1' after 282991200 ps,
'0' after 283073200 ps,
'1' after 283153200 ps,
'0' after 283236 ns,
'1' after 283315200 ps,
'0' after 283398400 ps,
'1' after 283478800 ps,
'0' after 283561600 ps,
'1' after 283640400 ps,
'0' after 283724 ns,
'1' after 283804400 ps,
'0' after 283887600 ps,
'1' after 283966 ns,
'0' after 284048800 ps,
'1' after 284130 ns,
'0' after 284212800 ps,
'1' after 284291200 ps,
'0' after 284374400 ps,
'1' after 284454800 ps,
'0' after 284538400 ps,
'1' after 284616800 ps,
'0' after 284699600 ps,
'1' after 284862400 ps,
'0' after 284945600 ps,
'1' after 285268400 ps,
'0' after 286166400 ps,
'1' after 286570400 ps,
'0' after 286980400 ps,
'1' after 287384800 ps,
'0' after 287794400 ps,
'1' after 288117600 ps,
'0' after 288200 ns,
'1' after 288443200 ps,
'0' after 288525600 ps,
'1' after 288606400 ps,
'0' after 288770400 ps,
'1' after 288849600 ps,
'0' after 288932800 ps,
'1' after 289012800 ps,
'0' after 289421600 ps,
'1' after 289825600 ps,
'0' after 290235600 ps,
'1' after 290640 ns,
'0' after 290967200 ps,
'1' after 291046800 ps,
'0' after 291212 ns,
'1' after 291372400 ps,
'0' after 291454800 ps,
'1' after 291535600 ps,
'0' after 291618800 ps,
'1' after 291697600 ps,
'0' after 291780800 ps,
'1' after 291860800 ps,
'0' after 291944400 ps,
'1' after 292022400 ps,
'0' after 292106 ns,
'1' after 292186800 ps,
'0' after 292269600 ps,
'1' after 292348 ns,
'0' after 292431600 ps,
'1' after 292512 ns,
'0' after 292595200 ps,
'1' after 292673600 ps,
'0' after 292756800 ps,
'1' after 292838 ns,
'0' after 292920400 ps,
'1' after 292999200 ps,
'0' after 293082800 ps,
'1' after 293162800 ps,
'0' after 293246400 ps,
'1' after 293324400 ps,
'0' after 293408 ns,
'1' after 293488400 ps,
'0' after 293571600 ps,
'1' after 293650400 ps,
'0' after 293897200 ps,
'1' after 293976 ns,
'0' after 294059200 ps,
'1' after 294138400 ps,
'0' after 294223200 ps,
'1' after 294300400 ps,
'0' after 294384800 ps,
'1' after 294465200 ps,
'0' after 294548400 ps,
'1' after 294626400 ps,
'0' after 294710 ns,
'1' after 294790400 ps,
'0' after 294873600 ps,
'1' after 294952400 ps,
'0' after 295035600 ps,
'1' after 295116 ns,
'0' after 295199200 ps,
'1' after 295277600 ps,
'0' after 295360800 ps,
'1' after 295442 ns,
'0' after 295524400 ps,
'1' after 295603200 ps,
'0' after 295768400 ps,
'1' after 295847600 ps,
'0' after 295930800 ps,
'1' after 296092 ns,
'0' after 296338 ns,
'1' after 296742400 ps,
'0' after 297151600 ps,
'1' after 297556 ns,
'0' after 297965200 ps,
'1' after 298207600 ps,
'0' after 298372400 ps,
'1' after 298452 ns,
'0' after 298616800 ps,
'1' after 298776800 ps,
'0' after 298859600 ps,
'1' after 298940400 ps,
'0' after 299023600 ps,
'1' after 299102400 ps,
'0' after 299184800 ps,
'1' after 299265600 ps,
'0' after 299348800 ps,
'1' after 299427600 ps,
'0' after 299510400 ps,
'1' after 299591200 ps,
'0' after 299674400 ps,
'1' after 299752800 ps,
'0' after 299836 ns,
'1' after 299916400 ps,
'0' after 300 us,
'1' after 300078400 ps,
'0' after 300161200 ps,
'1' after 300241600 ps,
'0' after 300325600 ps,
'1' after 300404 ns,
'0' after 300486800 ps,
'1' after 300567600 ps,
'0' after 300732 ns,
'1' after 300811200 ps,
'0' after 300894400 ps,
'1' after 300974400 ps,
'0' after 301139200 ps,
'1' after 301217600 ps,
'0' after 301300800 ps,
'1' after 301381600 ps,
'0' after 301464400 ps,
'1' after 301543200 ps,
'0' after 301626 ns,
'1' after 301706400 ps,
'0' after 301706800 ps,
'1' after 301707200 ps,
'0' after 301790 ns,
'1' after 301869200 ps,
'0' after 301952 ns,
'1' after 302032 ns,
'0' after 302115200 ps,
'1' after 302194400 ps,
'0' after 302276800 ps,
'1' after 302358 ns,
'0' after 302440800 ps,
'1' after 302519600 ps,
'0' after 302602800 ps,
'1' after 302683200 ps,
'0' after 302766400 ps,
'1' after 302845600 ps,
'0' after 302928 ns,
'1' after 303090 ns,
'0' after 303174 ns,
'1' after 303251600 ps,
'0' after 303416800 ps,
'1' after 303496800 ps,
'0' after 303661600 ps,
'1' after 304065600 ps,
'0' after 304475600 ps,
'1' after 304879200 ps,
'0' after 305289200 ps,
'1' after 305530800 ps,
'0' after 305695200 ps,
'1' after 305774800 ps,
'0' after 305775200 ps,
'1' after 305775600 ps,
'0' after 305940 ns,
'1' after 306018800 ps,
'0' after 306102400 ps,
'1' after 306994800 ps,
'0' after 307405600 ps,
'1' after 307484800 ps,
'0' after 307567200 ps,
'1' after 307647600 ps,
'0' after 307731200 ps,
'1' after 307809600 ps,
'0' after 307892400 ps,
'1' after 307973600 ps,
'0' after 308056400 ps,
'1' after 308135200 ps,
'0' after 308218 ns,
'1' after 308298800 ps,
'0' after 308382400 ps,
'1' after 308461200 ps,
'0' after 308544 ns,
'1' after 308624800 ps,
'0' after 308707600 ps,
'1' after 308786800 ps,
'0' after 308869600 ps,
'1' after 308949600 ps,
'0' after 309034 ns,
'1' after 309112400 ps,
'0' after 309276800 ps,
'1' after 309438400 ps,
'0' after 309684 ns,
'1' after 309844800 ps,
'0' after 309927600 ps,
'1' after 310008 ns,
'0' after 310091200 ps,
'1' after 310170 ns,
'0' after 310252800 ps,
'1' after 310333200 ps,
'0' after 310416800 ps,
'1' after 310494400 ps,
'0' after 310578 ns,
'1' after 310658800 ps,
'0' after 310742 ns,
'1' after 310821200 ps,
'0' after 310904400 ps,
'1' after 310984400 ps,
'0' after 311068400 ps,
'1' after 311145600 ps,
'0' after 311229600 ps,
'1' after 311310400 ps,
'0' after 311393200 ps,
'1' after 311472 ns,
'0' after 311554800 ps,
'1' after 311635200 ps,
'0' after 311718800 ps,
'1' after 311878800 ps,
'0' after 312043600 ps,
'1' after 312204800 ps,
'0' after 312287200 ps,
'1' after 312367600 ps,
'0' after 312450800 ps,
'1' after 312529200 ps,
'0' after 312612800 ps,
'1' after 312693600 ps,
'0' after 312776400 ps,
'1' after 312855200 ps,
'0' after 312938 ns,
'1' after 313018800 ps,
'0' after 313102400 ps,
'1' after 313180400 ps,
'0' after 313264 ns,
'1' after 313344 ns,
'0' after 313427200 ps,
'1' after 313505200 ps,
'0' after 313588800 ps,
'1' after 313670 ns,
'0' after 313752800 ps,
'1' after 313831200 ps,
'0' after 313914400 ps,
'1' after 314076800 ps,
'0' after 314160 ns,
'1' after 314238400 ps,
'0' after 314320800 ps,
'1' after 314402400 ps,
'0' after 314484800 ps,
'1' after 314564400 ps,
'0' after 314729200 ps,
'1' after 314808400 ps,
'0' after 314892 ns,
'1' after 314970800 ps,
'0' after 315054400 ps,
'1' after 315133200 ps,
'0' after 315216400 ps,
'1' after 315296400 ps,
'0' after 315380400 ps,
'1' after 315458800 ps,
'0' after 315542 ns,
'1' after 315622400 ps,
'0' after 315622800 ps,
'1' after 315623200 ps,
'0' after 315705600 ps,
'1' after 315784 ns,
'0' after 315867600 ps,
'1' after 315948 ns,
'0' after 316031200 ps,
'1' after 316109600 ps,
'0' after 316192800 ps,
'1' after 316273200 ps,
'0' after 316356400 ps,
'1' after 316435200 ps,
'0' after 316682 ns,
'1' after 316760800 ps,
'0' after 316844400 ps,
'1' after 317005600 ps,
'0' after 317170400 ps,
'1' after 317249200 ps,
'0' after 317332800 ps,
'1' after 317412400 ps,
'0' after 317496400 ps,
'1' after 317574 ns,
'0' after 317656800 ps,
'1' after 317738 ns,
'0' after 317821200 ps,
'1' after 317900 ns,
'0' after 317982800 ps,
'1' after 318063600 ps,
'0' after 318146800 ps,
'1' after 318225600 ps,
'0' after 318308400 ps,
'1' after 318389200 ps,
'0' after 318472400 ps,
'1' after 318550800 ps,
'0' after 318634400 ps,
'1' after 318714400 ps,
'0' after 318798 ns,
'1' after 318876 ns,
'0' after 318959600 ps,
'1' after 319040 ns,
'0' after 319123600 ps,
'1' after 319202 ns,
'0' after 319284800 ps,
'1' after 319447600 ps,
'0' after 319611600 ps,
'1' after 319690400 ps,
'0' after 319773200 ps,
'1' after 319853600 ps,
'0' after 319937200 ps,
'1' after 320015200 ps,
'0' after 320098400 ps,
'1' after 320179200 ps,
'0' after 320262 ns,
'1' after 320341200 ps,
'0' after 320424 ns,
'1' after 320504400 ps,
'0' after 320588400 ps,
'1' after 320666 ns,
'0' after 320749600 ps,
'1' after 320830400 ps,
'0' after 320913200 ps,
'1' after 320992 ns,
'0' after 321075200 ps,
'1' after 321155200 ps,
'0' after 321238800 ps,
'1' after 321317200 ps,
'0' after 321317600 ps,
'1' after 321318 ns,
'0' after 321482800 ps,
'1' after 321562400 ps,
'0' after 321645600 ps,
'1' after 321724 ns,
'0' after 321889200 ps,
'1' after 321968800 ps,
'0' after 322053600 ps,
'1' after 322456 ns,
'0' after 322866400 ps,
'1' after 323270 ns,
'0' after 323679600 ps,
'1' after 323840800 ps,
'0' after 324087200 ps,
'1' after 324247200 ps,
'0' after 324329200 ps,
'1' after 324492800 ps,
'0' after 324900400 ps,
'1' after 325304800 ps,
'0' after 325714800 ps,
'1' after 326118400 ps,
'0' after 326528 ns,
'1' after 326932800 ps,
'0' after 327830800 ps,
'1' after 328234800 ps,
'0' after 328644800 ps,
'1' after 329049200 ps,
'0' after 329458800 ps,
'1' after 329862 ns,
'0' after 330028 ns,
'1' after 330106400 ps,
'0' after 330272 ns,
'1' after 330350800 ps,
'0' after 330434800 ps,
'1' after 330676800 ps,
'0' after 331086400 ps,
'1' after 331490 ns,
'0' after 331899600 ps,
'1' after 332304 ns,
'0' after 332387200 ps,
'1' after 332712 ns,
'0' after 332875600 ps,
'1' after 333038 ns,
'0' after 333120400 ps,
'1' after 333524 ns,
'0' after 333933600 ps,
'1' after 334338400 ps,
'0' after 334748 ns,
'1' after 334989600 ps,
'0' after 335154400 ps,
'1' after 335233600 ps,
'0' after 335398800 ps,
'1' after 335559600 ps,
'0' after 335968 ns,
'1' after 336372400 ps,
'0' after 336781600 ps,
'1' after 337186 ns,
'0' after 337268800 ps,
'1' after 337349600 ps,
'0' after 337514 ns,
'1' after 337593200 ps,
'0' after 337676400 ps,
'1' after 337838 ns,
'0' after 338002400 ps,
'1' after 338081200 ps,
'0' after 338164800 ps,
'1' after 338244 ns,
'0' after 338327200 ps,
'1' after 338407200 ps,
'0' after 338490800 ps,
'1' after 338569200 ps,
'0' after 338652400 ps,
'1' after 338733200 ps,
'0' after 338816 ns,
'1' after 338895200 ps,
'0' after 338978400 ps,
'1' after 339058400 ps,
'0' after 339142 ns,
'1' after 339219600 ps,
'0' after 339303600 ps,
'1' after 339384400 ps,
'0' after 339467200 ps,
'1' after 339546400 ps,
'0' after 339629200 ps,
'1' after 339709600 ps,
'0' after 339793200 ps,
'1' after 339952400 ps,
'0' after 340035600 ps,
'1' after 340116400 ps,
'0' after 340362400 ps,
'1' after 340441200 ps,
'0' after 340525600 ps,
'1' after 340602400 ps,
'0' after 340602800 ps,
'1' after 340603200 ps,
'0' after 340686400 ps,
'1' after 340767600 ps,
'0' after 340850 ns,
'1' after 340929600 ps,
'0' after 341012400 ps,
'1' after 341092800 ps,
'0' after 341176400 ps,
'1' after 341254400 ps,
'0' after 341338 ns,
'1' after 341418 ns,
'0' after 341501200 ps,
'1' after 341580 ns,
'0' after 341663200 ps,
'1' after 341743600 ps,
'0' after 341827200 ps,
'1' after 341905600 ps,
'0' after 341988800 ps,
'1' after 342069200 ps,
'0' after 342152400 ps,
'1' after 342230800 ps,
'0' after 342314 ns,
'1' after 342395200 ps,
'0' after 342478 ns,
'1' after 342557200 ps,
'0' after 342639600 ps,
'1' after 342801600 ps,
'0' after 342885200 ps,
'1' after 342963200 ps,
'0' after 343046 ns,
'1' after 343127200 ps,
'0' after 343210 ns,
'1' after 343288800 ps,
'0' after 343372 ns,
'1' after 343452 ns,
'0' after 343536 ns,
'1' after 343614400 ps,
'0' after 343697200 ps,
'1' after 343777600 ps,
'0' after 343861200 ps,
'1' after 343940 ns,
'0' after 344022800 ps,
'1' after 344104 ns,
'0' after 344186800 ps,
'1' after 344265200 ps,
'0' after 344348800 ps,
'1' after 344428800 ps,
'0' after 344512400 ps,
'1' after 344590400 ps,
'0' after 344673600 ps,
'1' after 344754400 ps,
'0' after 344919200 ps,
'1' after 345323200 ps,
'0' after 345323600 ps,
'1' after 345324 ns,
'0' after 345732800 ps,
'1' after 346137200 ps,
'0' after 346546400 ps,
'1' after 346950400 ps,
'0' after 347360 ns,
'1' after 347438800 ps,
'0' after 347523200 ps,
'1' after 347601600 ps,
'0' after 347684400 ps,
'1' after 347765600 ps,
'0' after 348662400 ps,
'1' after 349066800 ps,
'0' after 349476800 ps,
'1' after 349881200 ps,
'0' after 350290800 ps,
'1' after 350694800 ps,
'0' after 350941600 ps,
'1' after 351020 ns,
'0' after 351104400 ps,
'1' after 351183200 ps,
'0' after 351430 ns,
'1' after 351508400 ps,
'0' after 351592800 ps,
'1' after 351671200 ps,
'0' after 351754800 ps,
'1' after 351834800 ps,
'0' after 351918800 ps,
'1' after 351996 ns,
'0' after 352079600 ps,
'1' after 352160400 ps,
'0' after 352243200 ps,
'1' after 352322400 ps,
'0' after 352405200 ps,
'1' after 352485600 ps,
'0' after 352568800 ps,
'1' after 352647200 ps,
'0' after 352730800 ps,
'1' after 352811600 ps,
'0' after 352894400 ps,
'1' after 352973200 ps,
'0' after 353056400 ps,
'1' after 353137200 ps,
'0' after 353383200 ps,
'1' after 353461600 ps,
'0' after 353544400 ps,
'1' after 353706400 ps,
'0' after 353871200 ps,
'1' after 353949600 ps,
'0' after 354033200 ps,
'1' after 354113200 ps,
'0' after 354196800 ps,
'1' after 354274800 ps,
'0' after 354358400 ps,
'1' after 354439600 ps,
'0' after 354522 ns,
'1' after 354600800 ps,
'0' after 354684 ns,
'1' after 354764400 ps,
'0' after 354847600 ps,
'1' after 354926 ns,
'0' after 355009200 ps,
'1' after 355090 ns,
'0' after 355172800 ps,
'1' after 355251600 ps,
'0' after 355334800 ps,
'1' after 355414800 ps,
'0' after 355498800 ps,
'1' after 355577200 ps,
'0' after 355660 ns,
'1' after 355984800 ps,
'0' after 356066800 ps,
'1' after 356148 ns,
'0' after 356393200 ps,
'1' after 356798 ns,
'0' after 357207200 ps,
'1' after 357611600 ps,
'0' after 358020800 ps,
'1' after 358181600 ps,
'0' after 358264400 ps,
'1' after 358344400 ps,
'0' after 358428 ns,
'1' after 358506400 ps,
'0' after 358589600 ps,
'1' after 358670800 ps,
'0' after 358834800 ps,
'1' after 359238800 ps,
'0' after 359648800 ps,
'1' after 360052800 ps,
'0' after 360462 ns,
'1' after 360622400 ps,
'0' after 360704800 ps,
'1' after 360868 ns,
'0' after 360950400 ps,
'1' after 361110800 ps,
'0' after 361274800 ps,
'1' after 361680800 ps,
'0' after 362089600 ps,
'1' after 362494 ns,
'0' after 362902800 ps,
'1' after 363144800 ps,
'0' after 363309600 ps,
'1' after 363389600 ps,
'0' after 363473200 ps,
'1' after 363551200 ps,
'0' after 363716400 ps,
'1' after 363796 ns,
'0' after 363880 ns,
'1' after 363957600 ps,
'0' after 363958 ns,
'1' after 363958400 ps,
'0' after 364041600 ps,
'1' after 364122400 ps,
'0' after 364204800 ps,
'1' after 364283600 ps,
'0' after 364367200 ps,
'1' after 364447600 ps,
'0' after 364530400 ps,
'1' after 364609600 ps,
'0' after 364692 ns,
'1' after 364773200 ps,
'0' after 364856 ns,
'1' after 364934800 ps,
'0' after 365018 ns,
'1' after 365098800 ps,
'0' after 365181200 ps,
'1' after 365260 ns,
'0' after 365343600 ps,
'1' after 365424400 ps,
'0' after 365507200 ps,
'1' after 365667600 ps,
'0' after 365750 ns,
'1' after 365830800 ps,
'0' after 365914 ns,
'1' after 365993200 ps,
'0' after 366158 ns,
'1' after 366237200 ps,
'0' after 366320400 ps,
'1' after 366399600 ps,
'0' after 366483600 ps,
'1' after 366561200 ps,
'0' after 366645200 ps,
'1' after 366726400 ps,
'0' after 366808800 ps,
'1' after 366887600 ps,
'0' after 366971200 ps,
'1' after 367051200 ps,
'0' after 367135200 ps,
'1' after 367212800 ps,
'0' after 367295600 ps,
'1' after 367376800 ps,
'0' after 367459200 ps,
'1' after 367538400 ps,
'0' after 367623600 ps,
'1' after 367701600 ps,
'0' after 367784400 ps,
'1' after 367864800 ps,
'0' after 367948400 ps,
'1' after 368027200 ps,
'0' after 368192 ns,
'1' after 368271200 ps,
'0' after 368355600 ps,
'1' after 368596400 ps,
'0' after 369494800 ps,
'1' after 369899200 ps,
'0' after 370309200 ps,
'1' after 370713600 ps,
'0' after 371122400 ps,
'1' after 371527200 ps,
'0' after 371936400 ps,
'1' after 372097200 ps,
'0' after 372179600 ps,
'1' after 372260 ns,
'0' after 372343200 ps,
'1' after 372421600 ps,
'0' after 372505600 ps,
'1' after 372585200 ps,
'0' after 372669200 ps,
'1' after 372747200 ps,
'0' after 372830400 ps,
'1' after 372911200 ps,
'0' after 372994 ns,
'1' after 373073200 ps,
'0' after 373156400 ps,
'1' after 373236 ns,
'0' after 373320 ns,
'1' after 373397600 ps,
'0' after 373481600 ps,
'1' after 373562400 ps,
'0' after 373645200 ps,
'1' after 373723600 ps,
'0' after 373806800 ps,
'1' after 373888 ns,
'0' after 373970800 ps,
'1' after 374049600 ps,
'0' after 374296 ns,
'1' after 374375200 ps,
'0' after 374459600 ps,
'1' after 374618800 ps,
'0' after 374701600 ps,
'1' after 374783200 ps,
'0' after 374865600 ps,
'1' after 374944400 ps,
'0' after 375028400 ps,
'1' after 375107200 ps,
'0' after 375190800 ps,
'1' after 375270800 ps,
'0' after 375354400 ps,
'1' after 375432400 ps,
'0' after 375516 ns,
'1' after 375596800 ps,
'0' after 375679200 ps,
'1' after 375758 ns,
'0' after 375841600 ps,
'1' after 375921600 ps,
'0' after 376005200 ps,
'1' after 376083200 ps,
'0' after 376166800 ps,
'1' after 376247600 ps,
'0' after 376330400 ps,
'1' after 376409200 ps,
'0' after 376492800 ps,
'1' after 376572800 ps,
'0' after 376818800 ps,
'1' after 377142 ns,
'0' after 377224400 ps,
'1' after 377630400 ps,
'0' after 378039200 ps,
'1' after 378443600 ps,
'0' after 378853200 ps,
'1' after 379257200 ps,
'0' after 379340 ns,
'1' after 379502800 ps,
'0' after 379585600 ps,
'1' after 379663600 ps,
'0' after 380074 ns,
'1' after 380477600 ps,
'0' after 380886800 ps,
'1' after 381291600 ps,
'0' after 381374400 ps,
'1' after 381618400 ps,
'0' after 381699600 ps,
'1' after 381944 ns,
'0' after 382025600 ps,
'1' after 382105600 ps,
'0' after 382514800 ps,
'1' after 382918400 ps,
'0' after 383328400 ps,
'1' after 383732800 ps,
'0' after 384060800 ps,
'1' after 384139600 ps,
'0' after 384386 ns,
'1' after 384546400 ps,
'0' after 384629600 ps,
'1' after 384709600 ps,
'0' after 384793200 ps,
'1' after 384871600 ps,
'0' after 384954800 ps,
'1' after 385035600 ps,
'0' after 385118400 ps,
'1' after 385197200 ps,
'0' after 385280400 ps,
'1' after 385361200 ps,
'0' after 385444 ns,
'1' after 385522400 ps,
'0' after 385606 ns,
'1' after 385686400 ps,
'0' after 385769600 ps,
'1' after 385848 ns,
'0' after 385931200 ps,
'1' after 386012 ns,
'0' after 386094800 ps,
'1' after 386174 ns,
'0' after 386256800 ps,
'1' after 386337600 ps,
'0' after 386420800 ps,
'1' after 386498800 ps,
'0' after 386582400 ps,
'1' after 386744400 ps,
'0' after 386828 ns,
'1' after 386987200 ps,
'0' after 387070 ns,
'1' after 387151600 ps,
'0' after 387234 ns,
'1' after 387313200 ps,
'0' after 387396400 ps,
'1' after 387476400 ps,
'0' after 387560400 ps,
'1' after 387638400 ps,
'0' after 387721200 ps,
'1' after 387802800 ps,
'0' after 387885200 ps,
'1' after 387964 ns,
'0' after 388047200 ps,
'1' after 388127600 ps,
'0' after 388211200 ps,
'1' after 388289600 ps,
'0' after 388372400 ps,
'1' after 388453600 ps,
'0' after 388536400 ps,
'1' after 388614800 ps,
'0' after 388698 ns,
'1' after 388778800 ps,
'0' after 388861600 ps,
'1' after 389022 ns,
'0' after 389186800 ps,
'1' after 389266400 ps,
'0' after 389350400 ps,
'1' after 389428400 ps,
'0' after 390326800 ps,
'1' after 390730400 ps,
'0' after 390814 ns,
'1' after 390895200 ps,
'0' after 390978 ns,
'1' after 391056800 ps,
'0' after 391140 ns,
'1' after 391220800 ps,
'0' after 391303600 ps,
'1' after 391382800 ps,
'0' after 391466 ns,
'1' after 391546 ns,
'0' after 391629200 ps,
'1' after 391708 ns,
'0' after 391791200 ps,
'1' after 391872 ns,
'0' after 391954800 ps,
'1' after 392033200 ps,
'0' after 392116800 ps,
'1' after 392197200 ps,
'0' after 392280 ns,
'1' after 392358800 ps,
'0' after 392524 ns,
'1' after 392603200 ps,
'0' after 392768800 ps,
'1' after 393010800 ps,
'0' after 393092800 ps,
'1' after 393174 ns,
'0' after 393582400 ps,
'1' after 393986800 ps,
'0' after 394396 ns,
'1' after 394799600 ps,
'0' after 395128400 ps,
'1' after 395207600 ps,
'0' after 395292 ns,
'1' after 395614 ns,
'0' after 396024 ns,
'1' after 396427600 ps,
'0' after 396837200 ps,
'1' after 397241600 ps,
'0' after 397406400 ps,
'1' after 397486 ns,
'0' after 397570 ns,
'1' after 397648 ns,
'0' after 398058 ns,
'1' after 398136 ns,
'0' after 398220 ns,
'1' after 398299200 ps,
'0' after 398383200 ps,
'1' after 398461200 ps,
'0' after 398544400 ps,
'1' after 398626 ns,
'0' after 398708 ns,
'1' after 398787200 ps,
'0' after 398870400 ps,
'1' after 398950800 ps,
'0' after 399034400 ps,
'1' after 399112400 ps,
'0' after 399196 ns,
'1' after 399276400 ps,
'0' after 399359600 ps,
'1' after 399438400 ps,
'0' after 399521600 ps,
'1' after 399602400 ps,
'0' after 399685200 ps,
'1' after 399764 ns,
'0' after 399847600 ps,
'1' after 399927200 ps;


		Instanz: ADAT_Taktgewinnung PORT MAP(clk => tb_clk,
														 In_ADAT => tb_Adat(0),
														 Out_ADAT_Clock => tb_AdatTakt,
														 Frame_Sync => tb_AdatFramesync
														 );
											
		C1: ADAT_Dekoder 
			generic map (AdatSchnittstellen => SCHNITTSTELLEN)
			PORT MAP(ADAT_Takt=> tb_AdatTakt,
						ADAT_Sync => to_bit(tb_AdatFramesync),
						In_ADAT => tb_adat,
						Out_Daten => tb_Out_Daten,
						Out_FrameOK => tb_Out_FrameOK
						);
  END;
